** Profile: "SCHEMATIC1-Bode1"  [ C:\Users\user\OneDrive\Desktop\Liron\Studies\PSPICE\PspiceAmplifierProject\PSPICE\amplifier-SCHEMATIC1-Bode1.sim ] 

** Creating circuit file "amplifier-SCHEMATIC1-Bode1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 0 1000
.PROBE 
.INC "../SCHEMATIC1.net"



.END
