** Profile: "SCHEMATIC1-Bode5"  [ C:\Users\user\OneDrive\Desktop\Liron\Studies\PSPICE\PspiceAmplifierProject\PSPICE\amplifier-SCHEMATIC1-Bode5.sim ] 

** Creating circuit file "amplifier-SCHEMATIC1-Bode5.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 1 10000
.PROBE 
.INC "amplifier-SCHEMATIC1.net" 

.INC "amplifier-SCHEMATIC1.als"


.END
