** Profile: "SCHEMATIC1-Bode6"  [ C:\Users\user\OneDrive\Desktop\Liron\Studies\PSPICE\PspiceAmplifierProject\PSPICE\amplifier-SCHEMATIC1-Bode6.sim ] 

** Creating circuit file "amplifier-SCHEMATIC1-Bode6.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 11 0.1 10000
.PROBE 
.INC "../SCHEMATIC1.net"



.END
