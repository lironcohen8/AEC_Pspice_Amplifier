** Profile: "SCHEMATIC1-sim1"  [ C:\Users\user\OneDrive\Desktop\Liron\Studies\PSPICE\amplifier-SCHEMATIC1-sim1.sim ] 

** Creating circuit file "amplifier-SCHEMATIC1-sim1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE 
.INC "../SCHEMATIC1.net"



.END
